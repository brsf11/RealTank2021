module Printer(input wire clk,rst_n,
               input wire);

endmodule