module NumShiftReg(input wire clk,rst_n,
                   input wire );

endmodule