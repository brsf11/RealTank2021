module Tube(input wire );

endmodule