module Printer();

endmodule